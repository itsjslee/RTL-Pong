module ball(
    input wire clk,
    output reg ball_direction
);

endmodule