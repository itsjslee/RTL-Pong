/* 
 * Pong Game Module
 * -------------------
 * This module controls the overall game logic
 * It handles:
 * - All modules
 */

module game (
    
)



