/* 
 * Pong Ball Module
 * -------------------
 * This module controls the ball movement in our Pong game.
 * It handles:
 * - Ball position tracking (x,y coordinates)
 * - Ball movement and direction
 * - Collision detection with paddles
 * - Screen boundary detection
 * - Reset functionality
 */

module ball
    input wire clk,
    input wire reset,
    output reg ball_direction
 

endmodule