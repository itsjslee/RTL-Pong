/* 
 * Pong Paddle Module
 * -------------------
 * This module controls the paddle movement in our Pong game.
 * It handles:
 * - Paddle position tracking (y coordinate)
 * - Paddle movement based on user input
 * - Screen boundary detection
 * - Reset functionality
 */

module paddle(
    input wire clk,
    input wire rst,
    input wire move_up,
    input wire move_down,
);

endmodule
